module orvl(x,y,z);
input x,y;
output z;
or g1(z,x,y);
endmodule