module xorvl(x,y,z);
input x,y;
output z;
xor g1(z,y,x);
endmodule