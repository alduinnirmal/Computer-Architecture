module andvl(x,y,z);
input x,y;
output z;
and g(z,y,x);
endmodule